module dff (
    input wire reset,
    input wire clk,
    input wire en,
    input wire d,
    output reg q
);

reg r_next, r_reg;

//memory part
always @ (posedge reset, posedge clk)
    begin 
        if (reset)
            r_reg <= 0;
        else 
            r_reg <= r_next;

    end

//next state logic
always @ (*)
    begin
        if (en) 
            r_next <= d;
        else 
            r_next <= r_reg;
    end

//output logic
always @ (*)
    begin
        q = r_reg;
    end


endmodule